`timescale 1ps/1ps

module s_box(
    input [3:0] x, 
    output [3:0] sx
    );

    assign sx[3] = (!x[3] & !x[1] & !x[0]) |
                   (!x[3] & x[1] & x[0]) |
                   (!x[3] & x[2] & !x[0]) |
                   (x[3] & !x[2] & x[0]) | 
                   (x[3] & !x[2] & x[1]);

    assign sx[2] = (!x[3] & !x[2] & !x[1]) | 
                   (!x[2] & !x[1] & x[0]) |
                   (!x[2] & x[1] & !x[0]) |
                   (x[3] & x[2] & !x[1]) |
                   (!x[3] & x[2] & x[1] & x[0]);
    
    assign sx[1] = (!x[3] & !x[2] & x[1]) | 
                   (!x[3] & x[1] & !x[0]) |
                   (!x[2] & x[1] & !x[0]) | 
                   (x[3] & !x[2] & !x[1]) |
                   (x[3] & x[2] & x[0]);

    assign sx[0] = (!x[3] & !x[2] & x[0]) |
                   (!x[3] & x[1] & x[0]) | 
                   (x[3] & !x[2] & !x[0]) |
                   (x[3] & x[2] & !x[0]) |
                   (!x[3] & x[2] & !x[1] & !x[0]) | 
                   (x[3] & x[2] & !x[1] & x[0]);

endmodule